../../../DAMIC/FPGA/ODILE_14/ethernet_firmware/top_ethernet.vhd